`timescale 10ns/100ps

module gamma_correction(
	input [6:0] red_in,
	input [6:0] green_in,
	input [5:0] blue_in,
	output reg [7:0] red_out,
	output reg [7:0] green_out,
	output reg [7:0] blue_out
);

always @(red_in) begin
	case (red_in)
		7'd0:	red_out = 8'd0;
		7'd1:	red_out = 8'd0;
		7'd2:	red_out = 8'd0;
		7'd3:	red_out = 8'd0;
		7'd4:	red_out = 8'd0;
		7'd5:	red_out = 8'd0;
		7'd6:	red_out = 8'd0;
		7'd7:	red_out = 8'd0;
		7'd8:	red_out = 8'd0;
		7'd9:	red_out = 8'd0;
		7'd10:	red_out = 8'd0;
		7'd11:	red_out = 8'd0;
		7'd12:	red_out = 8'd0;
		7'd13:	red_out = 8'd0;
		7'd14:	red_out = 8'd1;
		7'd15:	red_out = 8'd1;
		7'd16:	red_out = 8'd1;
		7'd17:	red_out = 8'd1;
		7'd18:	red_out = 8'd1;
		7'd19:	red_out = 8'd1;
		7'd20:	red_out = 8'd1;
		7'd21:	red_out = 8'd2;
		7'd22:	red_out = 8'd2;
		7'd23:	red_out = 8'd2;
		7'd24:	red_out = 8'd2;
		7'd25:	red_out = 8'd3;
		7'd26:	red_out = 8'd3;
		7'd27:	red_out = 8'd3;
		7'd28:	red_out = 8'd4;
		7'd29:	red_out = 8'd4;
		7'd30:	red_out = 8'd4;
		7'd31:	red_out = 8'd5;
		7'd32:	red_out = 8'd5;
		7'd33:	red_out = 8'd6;
		7'd34:	red_out = 8'd6;
		7'd35:	red_out = 8'd7;
		7'd36:	red_out = 8'd7;
		7'd37:	red_out = 8'd8;
		7'd38:	red_out = 8'd9;
		7'd39:	red_out = 8'd9;
		7'd40:	red_out = 8'd10;
		7'd41:	red_out = 8'd11;
		7'd42:	red_out = 8'd12;
		7'd43:	red_out = 8'd12;
		7'd44:	red_out = 8'd13;
		7'd45:	red_out = 8'd14;
		7'd46:	red_out = 8'd15;
		7'd47:	red_out = 8'd16;
		7'd48:	red_out = 8'd17;
		7'd49:	red_out = 8'd18;
		7'd50:	red_out = 8'd19;
		7'd51:	red_out = 8'd20;
		7'd52:	red_out = 8'd21;
		7'd53:	red_out = 8'd22;
		7'd54:	red_out = 8'd23;
		7'd55:	red_out = 8'd24;
		7'd56:	red_out = 8'd26;
		7'd57:	red_out = 8'd27;
		7'd58:	red_out = 8'd28;
		7'd59:	red_out = 8'd30;
		7'd60:	red_out = 8'd31;
		7'd61:	red_out = 8'd33;
		7'd62:	red_out = 8'd34;
		7'd63:	red_out = 8'd36;
		7'd64:	red_out = 8'd37;
		7'd65:	red_out = 8'd39;
		7'd66:	red_out = 8'd41;
		7'd67:	red_out = 8'd43;
		7'd68:	red_out = 8'd44;
		7'd69:	red_out = 8'd46;
		7'd70:	red_out = 8'd48;
		7'd71:	red_out = 8'd50;
		7'd72:	red_out = 8'd52;
		7'd73:	red_out = 8'd54;
		7'd74:	red_out = 8'd56;
		7'd75:	red_out = 8'd58;
		7'd76:	red_out = 8'd61;
		7'd77:	red_out = 8'd63;
		7'd78:	red_out = 8'd65;
		7'd79:	red_out = 8'd67;
		7'd80:	red_out = 8'd70;
		7'd81:	red_out = 8'd72;
		7'd82:	red_out = 8'd75;
		7'd83:	red_out = 8'd78;
		7'd84:	red_out = 8'd80;
		7'd85:	red_out = 8'd83;
		7'd86:	red_out = 8'd86;
		7'd87:	red_out = 8'd88;
		7'd88:	red_out = 8'd91;
		7'd89:	red_out = 8'd94;
		7'd90:	red_out = 8'd97;
		7'd91:	red_out = 8'd100;
		7'd92:	red_out = 8'd103;
		7'd93:	red_out = 8'd107;
		7'd94:	red_out = 8'd110;
		7'd95:	red_out = 8'd113;
		7'd96:	red_out = 8'd116;
		7'd97:	red_out = 8'd120;
		7'd98:	red_out = 8'd123;
		7'd99:	red_out = 8'd127;
		7'd100:	red_out = 8'd131;
		7'd101:	red_out = 8'd134;
		7'd102:	red_out = 8'd138;
		7'd103:	red_out = 8'd142;
		7'd104:	red_out = 8'd146;
		7'd105:	red_out = 8'd150;
		7'd106:	red_out = 8'd154;
		7'd107:	red_out = 8'd158;
		7'd108:	red_out = 8'd162;
		7'd109:	red_out = 8'd166;
		7'd110:	red_out = 8'd171;
		7'd111:	red_out = 8'd175;
		7'd112:	red_out = 8'd179;
		7'd113:	red_out = 8'd184;
		7'd114:	red_out = 8'd188;
		7'd115:	red_out = 8'd193;
		7'd116:	red_out = 8'd198;
		7'd117:	red_out = 8'd203;
		7'd118:	red_out = 8'd208;
		7'd119:	red_out = 8'd213;
		7'd120:	red_out = 8'd218;
		7'd121:	red_out = 8'd223;
		7'd122:	red_out = 8'd228;
		7'd123:	red_out = 8'd233;
		7'd124:	red_out = 8'd238;
		7'd125:	red_out = 8'd244;
		7'd126:	red_out = 8'd249;
		7'd127:	red_out = 8'd255;
	endcase
end


always @(green_in) begin
	case (green_in)
		7'd0:	green_out = 8'd0;
		7'd1:	green_out = 8'd0;
		7'd2:	green_out = 8'd0;
		7'd3:	green_out = 8'd0;
		7'd4:	green_out = 8'd0;
		7'd5:	green_out = 8'd0;
		7'd6:	green_out = 8'd0;
		7'd7:	green_out = 8'd0;
		7'd8:	green_out = 8'd0;
		7'd9:	green_out = 8'd0;
		7'd10:	green_out = 8'd0;
		7'd11:	green_out = 8'd0;
		7'd12:	green_out = 8'd0;
		7'd13:	green_out = 8'd0;
		7'd14:	green_out = 8'd1;
		7'd15:	green_out = 8'd1;
		7'd16:	green_out = 8'd1;
		7'd17:	green_out = 8'd1;
		7'd18:	green_out = 8'd1;
		7'd19:	green_out = 8'd1;
		7'd20:	green_out = 8'd1;
		7'd21:	green_out = 8'd2;
		7'd22:	green_out = 8'd2;
		7'd23:	green_out = 8'd2;
		7'd24:	green_out = 8'd2;
		7'd25:	green_out = 8'd3;
		7'd26:	green_out = 8'd3;
		7'd27:	green_out = 8'd3;
		7'd28:	green_out = 8'd4;
		7'd29:	green_out = 8'd4;
		7'd30:	green_out = 8'd4;
		7'd31:	green_out = 8'd5;
		7'd32:	green_out = 8'd5;
		7'd33:	green_out = 8'd6;
		7'd34:	green_out = 8'd6;
		7'd35:	green_out = 8'd7;
		7'd36:	green_out = 8'd7;
		7'd37:	green_out = 8'd8;
		7'd38:	green_out = 8'd9;
		7'd39:	green_out = 8'd9;
		7'd40:	green_out = 8'd10;
		7'd41:	green_out = 8'd11;
		7'd42:	green_out = 8'd12;
		7'd43:	green_out = 8'd12;
		7'd44:	green_out = 8'd13;
		7'd45:	green_out = 8'd14;
		7'd46:	green_out = 8'd15;
		7'd47:	green_out = 8'd16;
		7'd48:	green_out = 8'd17;
		7'd49:	green_out = 8'd18;
		7'd50:	green_out = 8'd19;
		7'd51:	green_out = 8'd20;
		7'd52:	green_out = 8'd21;
		7'd53:	green_out = 8'd22;
		7'd54:	green_out = 8'd23;
		7'd55:	green_out = 8'd24;
		7'd56:	green_out = 8'd26;
		7'd57:	green_out = 8'd27;
		7'd58:	green_out = 8'd28;
		7'd59:	green_out = 8'd30;
		7'd60:	green_out = 8'd31;
		7'd61:	green_out = 8'd33;
		7'd62:	green_out = 8'd34;
		7'd63:	green_out = 8'd36;
		7'd64:	green_out = 8'd37;
		7'd65:	green_out = 8'd39;
		7'd66:	green_out = 8'd41;
		7'd67:	green_out = 8'd43;
		7'd68:	green_out = 8'd44;
		7'd69:	green_out = 8'd46;
		7'd70:	green_out = 8'd48;
		7'd71:	green_out = 8'd50;
		7'd72:	green_out = 8'd52;
		7'd73:	green_out = 8'd54;
		7'd74:	green_out = 8'd56;
		7'd75:	green_out = 8'd58;
		7'd76:	green_out = 8'd61;
		7'd77:	green_out = 8'd63;
		7'd78:	green_out = 8'd65;
		7'd79:	green_out = 8'd67;
		7'd80:	green_out = 8'd70;
		7'd81:	green_out = 8'd72;
		7'd82:	green_out = 8'd75;
		7'd83:	green_out = 8'd78;
		7'd84:	green_out = 8'd80;
		7'd85:	green_out = 8'd83;
		7'd86:	green_out = 8'd86;
		7'd87:	green_out = 8'd88;
		7'd88:	green_out = 8'd91;
		7'd89:	green_out = 8'd94;
		7'd90:	green_out = 8'd97;
		7'd91:	green_out = 8'd100;
		7'd92:	green_out = 8'd103;
		7'd93:	green_out = 8'd107;
		7'd94:	green_out = 8'd110;
		7'd95:	green_out = 8'd113;
		7'd96:	green_out = 8'd116;
		7'd97:	green_out = 8'd120;
		7'd98:	green_out = 8'd123;
		7'd99:	green_out = 8'd127;
		7'd100:	green_out = 8'd131;
		7'd101:	green_out = 8'd134;
		7'd102:	green_out = 8'd138;
		7'd103:	green_out = 8'd142;
		7'd104:	green_out = 8'd146;
		7'd105:	green_out = 8'd150;
		7'd106:	green_out = 8'd154;
		7'd107:	green_out = 8'd158;
		7'd108:	green_out = 8'd162;
		7'd109:	green_out = 8'd166;
		7'd110:	green_out = 8'd171;
		7'd111:	green_out = 8'd175;
		7'd112:	green_out = 8'd179;
		7'd113:	green_out = 8'd184;
		7'd114:	green_out = 8'd188;
		7'd115:	green_out = 8'd193;
		7'd116:	green_out = 8'd198;
		7'd117:	green_out = 8'd203;
		7'd118:	green_out = 8'd208;
		7'd119:	green_out = 8'd213;
		7'd120:	green_out = 8'd218;
		7'd121:	green_out = 8'd223;
		7'd122:	green_out = 8'd228;
		7'd123:	green_out = 8'd233;
		7'd124:	green_out = 8'd238;
		7'd125:	green_out = 8'd244;
		7'd126:	green_out = 8'd249;
		7'd127:	green_out = 8'd255;
	endcase
end


always @(blue_in) begin
	case (blue_in)
		6'd0:	blue_out = 8'd0;
		6'd1:	blue_out = 8'd0;
		6'd2:	blue_out = 8'd0;
		6'd3:	blue_out = 8'd0;
		6'd4:	blue_out = 8'd0;
		6'd5:	blue_out = 8'd0;
		6'd6:	blue_out = 8'd0;
		6'd7:	blue_out = 8'd1;
		6'd8:	blue_out = 8'd1;
		6'd9:	blue_out = 8'd1;
		6'd10:	blue_out = 8'd1;
		6'd11:	blue_out = 8'd2;
		6'd12:	blue_out = 8'd2;
		6'd13:	blue_out = 8'd3;
		6'd14:	blue_out = 8'd4;
		6'd15:	blue_out = 8'd5;
		6'd16:	blue_out = 8'd5;
		6'd17:	blue_out = 8'd7;
		6'd18:	blue_out = 8'd8;
		6'd19:	blue_out = 8'd9;
		6'd20:	blue_out = 8'd10;
		6'd21:	blue_out = 8'd12;
		6'd22:	blue_out = 8'd13;
		6'd23:	blue_out = 8'd15;
		6'd24:	blue_out = 8'd17;
		6'd25:	blue_out = 8'd19;
		6'd26:	blue_out = 8'd21;
		6'd27:	blue_out = 8'd24;
		6'd28:	blue_out = 8'd26;
		6'd29:	blue_out = 8'd29;
		6'd30:	blue_out = 8'd32;
		6'd31:	blue_out = 8'd35;
		6'd32:	blue_out = 8'd38;
		6'd33:	blue_out = 8'd42;
		6'd34:	blue_out = 8'd45;
		6'd35:	blue_out = 8'd49;
		6'd36:	blue_out = 8'd53;
		6'd37:	blue_out = 8'd57;
		6'd38:	blue_out = 8'd62;
		6'd39:	blue_out = 8'd67;
		6'd40:	blue_out = 8'd71;
		6'd41:	blue_out = 8'd77;
		6'd42:	blue_out = 8'd82;
		6'd43:	blue_out = 8'd88;
		6'd44:	blue_out = 8'd93;
		6'd45:	blue_out = 8'd99;
		6'd46:	blue_out = 8'd106;
		6'd47:	blue_out = 8'd112;
		6'd48:	blue_out = 8'd119;
		6'd49:	blue_out = 8'd126;
		6'd50:	blue_out = 8'd134;
		6'd51:	blue_out = 8'd141;
		6'd52:	blue_out = 8'd149;
		6'd53:	blue_out = 8'd157;
		6'd54:	blue_out = 8'd166;
		6'd55:	blue_out = 8'd174;
		6'd56:	blue_out = 8'd183;
		6'd57:	blue_out = 8'd193;
		6'd58:	blue_out = 8'd202;
		6'd59:	blue_out = 8'd212;
		6'd60:	blue_out = 8'd222;
		6'd61:	blue_out = 8'd233;
		6'd62:	blue_out = 8'd244;
		6'd63:	blue_out = 8'd255;
	endcase
end

endmodule